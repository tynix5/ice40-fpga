module ps2_top(

);

endmodule