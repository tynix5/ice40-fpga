module main(input switch, output led);

assign led = switch;

endmodule