module pong_score(

    input [3:0] score,      // 0-9
    output [349:0] state    // 35x10 bitmap
);

    // digits 0-9 bitmap
    // size of original font 7x5 --> 7x10 due to half clock speed
    // size of each character on display increased to 35x10 (technically 35x25)
    reg [349:0] digit_bitmap[9:0];

    initial begin

        digit_bitmap[0] <= {{5{10'b0011111100}}, {5{10'b1100000011}}, {5{10'b1100001111}}, {5{10'b1100110011}}, {5{10'b1111000011}}, {5{10'b1100000011}}, {5{10'b0011111100}}};
        digit_bitmap[1] <= {{5{10'b1111111111}}, {5{10'b0000110000}}, {5{10'b0000110000}}, {5{10'b0000110000}}, {5{10'b0000110000}}, {5{10'b0000111100}}, {5{10'b0000110000}}};
        digit_bitmap[2] <= {{5{10'b1111111111}}, {5{10'b0000000011}}, {5{10'b0000001100}}, {5{10'b0011110000}}, {5{10'b1100000000}}, {5{10'b1100000011}}, {5{10'b0011111100}}};
        digit_bitmap[3] <= {{5{10'b0011111100}}, {5{10'b1100000011}}, {5{10'b1100000000}}, {5{10'b0011110000}}, {5{10'b0011000000}}, {5{10'b1100000000}}, {5{10'b1111111111}}};
        digit_bitmap[4] <= {{5{10'b0011000000}}, {5{10'b0011000000}}, {5{10'b1111111111}}, {5{10'b0011000011}}, {5{10'b0011001100}}, {5{10'b0011110000}}, {5{10'b0011000000}}};
        digit_bitmap[5] <= {{5{10'b0011111100}}, {5{10'b1100000011}}, {5{10'b1100000000}}, {5{10'b1100000000}}, {5{10'b0011111111}}, {5{10'b0000000011}}, {5{10'b1111111111}}};
        digit_bitmap[6] <= {{5{10'b0011111100}}, {5{10'b1100000011}}, {5{10'b1100000011}}, {5{10'b0011111111}}, {5{10'b0000000011}}, {5{10'b0000001100}}, {5{10'b1111110000}}};
        digit_bitmap[7] <= {{5{10'b0000001100}}, {5{10'b0000001100}}, {5{10'b0000001100}}, {5{10'b0000110000}}, {5{10'b0011000000}}, {5{10'b1100000000}}, {5{10'b1111111111}}};
        digit_bitmap[8] <= {{5{10'b0011111100}}, {5{10'b1100000011}}, {5{10'b1100000011}}, {5{10'b0011111100}}, {5{10'b1100000011}}, {5{10'b1100000011}}, {5{10'b0011111100}}};
        digit_bitmap[9] <= {{5{10'b0000111111}}, {5{10'b0011000000}}, {5{10'b1100000000}}, {5{10'b1111111100}}, {5{10'b1100000011}}, {5{10'b1100000011}}, {5{10'b0011111100}}};

    end

    assign state = (score < 10) ? digit_bitmap[score] : 350'b0;

endmodule