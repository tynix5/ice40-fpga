module pong_score(

    input clk,
    input rst,
    input [3:0] score,      // 0-9
    output [34:0] state
);

    // 10x7x5 score
    reg [34:0] score_mem[9:0];

    initial begin

        score_mem[0] <= 35'b01110100011001110101110011000101110;
        score_mem[1] <= 35'b01110001000010000100001000011000100;
        score_mem[2] <= 35'b11111000010001001100100001000101110;
        score_mem[3] <= 35'b01110100011000001100010001000011111;
        score_mem[4] <= 35'b01000010001111101001010100110001000;
        score_mem[5] <= 35'b01110100011000010000011110000111111;
        score_mem[6] <= 35'b01110100011000101111000010001011100;
        score_mem[7] <= 35'b00010000100001000100010001000011111;
        score_mem[8] <= 35'b01110100011000101110100011000101110;
        score_mem[9] <= 35'b00111010001000011110100011000101110;

    end

    assign state = (score < 10) ? score_mem[score] : 35'b0;

endmodule